../../../rtl/frame_generator/frame_generator_impl.sv