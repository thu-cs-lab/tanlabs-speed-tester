../../../rtl/tester_common.svh