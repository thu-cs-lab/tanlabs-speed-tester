../../../rtl/frame_checker/frame_checker_impl.sv